// ----------------------
// Instruction Decoder
// ----------------------
module instruction_decoder(
    input  [31:0] instruction,
    output reg [4:0]  opcode, 
    output reg [4:0]  rd,    
    output reg [4:0]  rs,    
    output reg [4:0]  rt,      
    output reg [11:0] literal, 
    output reg [3:0]  alu_op,
    output reg        is_immediate,
    output reg        reg_write_enable,
    output reg        is_float
);
    localparam ALU_ADD  = 4'b0000;
    localparam ALU_SUB  = 4'b0001;
    localparam ALU_MUL  = 4'b0010;
    localparam ALU_DIV  = 4'b0011;
    localparam ALU_SHR  = 4'b0100;
    localparam ALU_SHL  = 4'b0101;
    localparam ALU_AND  = 4'b0110;
    localparam ALU_OR   = 4'b0111;
    localparam ALU_XOR  = 4'b1000;
    localparam ALU_NOT  = 4'b1001;
    always @(*) begin
        opcode   = instruction[31:27];
        rd       = instruction[26:22];
        rs       = instruction[21:17];
        rt       = instruction[16:12];
        literal  = instruction[11:0];
        is_immediate     = 0;
        reg_write_enable = 1;
        is_float         = 0;
        alu_op           = ALU_ADD;
        case (opcode)
            5'b11000: alu_op = ALU_ADD;
            5'b11001: begin alu_op = ALU_ADD; is_immediate = 1; end
            5'b11010: alu_op = ALU_SUB;
            5'b11011: begin alu_op = ALU_SUB; is_immediate = 1; end
            5'b11100: alu_op = ALU_MUL;
            5'b11101: alu_op = ALU_DIV;
            5'b00000: alu_op = ALU_AND;
            5'b00001: alu_op = ALU_OR;
            5'b00010: alu_op = ALU_XOR;
            5'b00011: alu_op = ALU_NOT;
            5'b00100: alu_op = ALU_SHR;
            5'b00101: begin alu_op = ALU_SHR; is_immediate = 1; end
            5'b00110: alu_op = ALU_SHL;
            5'b00111: begin alu_op = ALU_SHL; is_immediate = 1; end
            5'b10001: begin alu_op = ALU_ADD; end
            5'b10010: begin alu_op = ALU_ADD; is_immediate = 1; end
            5'b10100: begin alu_op = ALU_ADD; is_float = 1; end
            5'b10101: begin alu_op = ALU_SUB; is_float = 1; end
            5'b10110: begin alu_op = ALU_MUL; is_float = 1; end
            5'b10111: begin alu_op = ALU_DIV; is_float = 1; end
            default: begin reg_write_enable = 0; end
        endcase
    end
endmodule

// ----------------------
// Register File
// ----------------------
module register_file(
    input clk,
    input  [4:0] rs_addr,
    input  [4:0] rt_addr,
    input  [4:0] rd_addr,
    input  [63:0] write_data,
    input         write_enable,
    output [63:0] rs_data,
    output [63:0] rt_data
);
    reg [63:0] registers [0:31];
    integer i;
    initial begin
        for (i = 0; i < 32; i = i + 1)
            registers[i] = 64'd0;
    end
    assign rs_data = registers[rs_addr];
    assign rt_data = registers[rt_addr];
    always @(posedge clk) begin
        if (write_enable && (rd_addr != 5'd0))
            registers[rd_addr] <= write_data;
    end
endmodule

// ----------------------
// Control Module
// ----------------------
module control(
    input [4:0] op,
    input [63:0] rd,
    input [63:0] rs,
    input [63:0] rt,
    input [63:0] lit,
    input [63:0] inputPc,
    input [63:0] memData,
    output reg [63:0] pc
);
    localparam BR = 5'b01000;
    localparam BRR_RD = 5'b01001;
    localparam BRR_L = 5'b01010;
    localparam BRNZ = 5'b01011;
    localparam CALL = 5'b01100;
    localparam RET = 5'b01101;
    localparam BRGT = 5'b01110;
    always @(*) begin
        case(op)
            BR:      pc = rd;
            BRR_RD:  pc = inputPc + rd;
            BRR_L:   pc = inputPc + $signed(lit);
            BRNZ:    pc = (rs != 0) ? rd : inputPc + 4;
            CALL:    pc = rd;
            RET:     pc = memData;
            BRGT:    pc = (rs > rt) ? rd : inputPc + 4;
            default: pc = inputPc + 4;
        endcase
    end
endmodule

// ----------------------
// ALU/FPU Combined
// ----------------------
module alu_fpu(
    input  [63:0] a,
    input  [63:0] b,
    input  [3:0]  op,
    input         is_float,
    output reg [63:0] result
);
    real float_a, float_b, float_res;
    localparam ALU_ADD = 4'b0000;
    localparam ALU_SUB = 4'b0001;
    localparam ALU_MUL = 4'b0010;
    localparam ALU_DIV = 4'b0011;
    localparam ALU_SHR = 4'b0100;
    localparam ALU_SHL = 4'b0101;
    localparam ALU_AND = 4'b0110;
    localparam ALU_OR  = 4'b0111;
    localparam ALU_XOR = 4'b1000;
    localparam ALU_NOT = 4'b1001;
    always @(*) begin
        if (is_float) begin
            float_a = $bitstoreal(a);
            float_b = $bitstoreal(b);
            case (op)
                ALU_ADD: float_res = float_a + float_b;
                ALU_SUB: float_res = float_a - float_b;
                ALU_MUL: float_res = float_a * float_b;
                ALU_DIV: float_res = float_a / float_b;
                default: float_res = 0.0;
            endcase
            result = $realtobits(float_res);
        end else begin
            case (op)
                ALU_ADD: result = a + b;
                ALU_SUB: result = a - b;
                ALU_MUL: result = a * b;
                ALU_DIV: result = (b != 0) ? (a / b) : 64'd0;
                ALU_SHR: result = a >> b[5:0];
                ALU_SHL: result = a << b[5:0];
                ALU_AND: result = a & b;
                ALU_OR : result = a | b;
                ALU_XOR: result = a ^ b;
                ALU_NOT: result = ~a;
                default: result = 64'd0;
            endcase
        end
    end
endmodule

// ----------------------
// Clock Generator
// ----------------------
module clock_generator(
    output reg clk
);
    initial begin
        clk = 0;
    end
    always begin
        #5 clk = ~clk;
    end
endmodule

// ----------------------
// Fetch Module
// ----------------------
module fetch(
    input clk,
    input reset,
    input [63:0] sp,
    input [63:0] new_pc,
    output reg [63:0] pc_out
);
    reg [63:0] curr_pc;
    assign pc_out = curr_pc;
    always @(posedge clk or posedge reset) begin
        if(reset)
            curr_pc <= 64'h2000;
        else
            curr_pc <= new_pc;
    end
endmodule

// ----------------------
// MemoryHandler Module
// ----------------------
module memoryHandler(
    input [4:0] opcode,
    input [63:0] rd, rs, lit, pc, r31,
    output reg [63:0] mem_addr,
    output reg [63:0] mem_wr_data,
    output reg mem_wr_en,
    output reg mem_reg_write
);
    always @(*) begin
        case(opcode)
            5'b01100: begin
                mem_addr = r31 - 8;
                mem_wr_data = pc + 4;
                mem_wr_en = 1;
                mem_reg_write = 0;
            end
            5'b01101: begin
                mem_addr = r31 - 8;
                mem_wr_data = 0;
                mem_wr_en = 0;
                mem_reg_write = 0;
            end
            5'b10000: begin
                mem_addr = rs + lit;
                mem_wr_data = 0;
                mem_wr_en = 0;
                mem_reg_write = 1;
            end
            5'b10011: begin
                mem_addr = rd + lit;
                mem_wr_data = rs;
                mem_wr_en = 1;
                mem_reg_write = 0;
            end
            default: begin
                mem_addr = 64'h2000;
                mem_wr_data = 0;
                mem_wr_en = 0;
                mem_reg_write = 0;
            end
        endcase
    end
endmodule

// ----------------------
// Memory Module
// ----------------------
module memory(
    input [63:0] addr_pc,
    input clk,
    input reset,
    input write_en,
    input [63:0] data_in,
    input [63:0] addr_rw,
    output reg [63:0] data_out,
    output reg [31:0] inst_out
);
    reg [7:0] bytes [0:524287];
    integer idx;
    always @(*) begin
        inst_out[7:0] = bytes[addr_pc];
        inst_out[15:8] = bytes[addr_pc+1];
        inst_out[23:16] = bytes[addr_pc+2];
        inst_out[31:24] = bytes[addr_pc+3];
    end
    always @(*) begin
        data_out[7:0] = bytes[addr_rw];
        data_out[15:8] = bytes[addr_rw+1];
        data_out[23:16] = bytes[addr_rw+2];
        data_out[31:24] = bytes[addr_rw+3];
        data_out[39:32] = bytes[addr_rw+4];
        data_out[47:40] = bytes[addr_rw+5];
        data_out[55:48] = bytes[addr_rw+6];
        data_out[63:56] = bytes[addr_rw+7];
    end
    always @(posedge clk or posedge reset) begin
        if(reset) begin
            for(idx = 0; idx < 524288; idx = idx + 1)
                bytes[idx] <= 8'b0;
        end else if(write_en) begin
            bytes[addr_rw] <= data_in[7:0];
            bytes[addr_rw+1] <= data_in[15:8];
            bytes[addr_rw+2] <= data_in[23:16];
            bytes[addr_rw+3] <= data_in[31:24];
            bytes[addr_rw+4] <= data_in[39:32];
            bytes[addr_rw+5] <= data_in[47:40];
            bytes[addr_rw+6] <= data_in[55:48];
            bytes[addr_rw+7] <= data_in[63:56];
        end
    end
endmodule

// ----------------------
// Reg-Literal Mux Module
// ----------------------
module reglitmux(
    input [4:0] sel,
    input [63:0] reg_val,
    input [63:0] imm_val,
    output reg [63:0] mux_out
);
    always @(*) begin
        case(sel)
            5'b11001, 5'b11011, 5'b00101, 5'b00111, 5'b10010: mux_out = imm_val;
            default: mux_out = reg_val;
        endcase
    end
endmodule

// ----------------------
// Top-Level Module: tinker_core
// ----------------------
module tinker_core(
    input clk,
    input reset
);
    wire [31:0] pc;
    wire branch = 1'b0;
    wire [31:0] branch_address = 32'd0;
    
    program_counter pc_inst(
        .clk(clk),
        .reset(reset),
        .branch(branch),
        .branch_address(branch_address),
        .pc(pc)
    );
    
    wire [31:0] instruction;
    instruction_fetch fetch_inst(
        .clk(clk),
        .reset(reset),
        .mem_read(1'b1),
        .instruction(instruction),
        .pc(pc)
    );
    
    wire [4:0] opcode, rd, rs, rt;
    wire [11:0] literal;
    wire [3:0] alu_op;
    wire is_immediate, reg_write_enable, is_float;
    instruction_decoder decoder_inst(
        .instruction(instruction),
        .opcode(opcode),
        .rd(rd),
        .rs(rs),
        .rt(rt),
        .literal(literal),
        .alu_op(alu_op),
        .is_immediate(is_immediate),
        .reg_write_enable(reg_write_enable),
        .is_float(is_float)
    );
    
    wire [63:0] rs_data, rt_data;
    register_file reg_file(
        .clk(clk),
        .rs_addr(rs),
        .rt_addr(rt),
        .rd_addr(rd),
        .write_data(result),
        .write_enable(reg_write_enable),
        .rs_data(rs_data),
        .rt_data(rt_data)
    );
    
    wire [63:0] result;
    wire [63:0] operand_b;
    assign operand_b = is_immediate ? {{52{literal[11]}}, literal} : rt_data;
    
    alu_fpu alu_unit(
        .a(rs_data),
        .b(operand_b),
        .op(alu_op),
        .is_float(is_float),
        .result(result)
    );
endmodule
